typedef uvm_sequencer #(fifo_rd_tx) fifo_rd_sequencer;
