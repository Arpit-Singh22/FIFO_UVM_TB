class fifo_common;
	static int wr_tx_count;
	static int wr_drv_count;
	static int matchings;
	static int mismatchings;
endclass
