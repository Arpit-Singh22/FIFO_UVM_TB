typedef uvm_sequencer #(fifo_wr_tx) fifo_wr_sequencer;
